library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MIPS is
    port (
        clk : in std_logic;
        reset : in std_logic;
    );
end MIPS;

architecture Behavioral of MIPS is
begin

end Behavioral;