library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ControlUnit is
    port (
        -- Inputs
        OP          : in  std_logic_vector(5 downto 0);  -- Opcode
        -- Funct input is removed
        
        -- Main Control Outputs
        RegWrite    : out std_logic;
        RegDst      : out std_logic;
        Branch      : out std_logic;
        MemRead     : out std_logic;
        MemtoReg    : out std_logic;
        MemWrite    : out std_logic;
        ALUSrc      : out std_logic;
        Jump        : out std_logic;
        
        -- Changed ALU Control Output to 2-bit ALUOp
        ALUOp_o     : out std_logic_vector(1 downto 0)
    );
end entity ControlUnit;

architecture Behavioral of ControlUnit is
    -- Internal signals
    signal ALUOp : std_logic_vector(1 downto 0); -- This signal is generated by the main control logic
begin
    -- Main Control Logic (determines ALUOp and other control signals)
    process(OP)
    begin
        case OP is
            -- R-type
            when "000000" =>
                RegWrite <= '1';
                RegDst   <= '1';
                Branch   <= '0';
                MemRead  <= '0';
                MemtoReg <= '0';
                MemWrite <= '0';
                ALUSrc   <= '0';
                Jump     <= '0';
                ALUOp    <= "10"; -- ALUOp for R-type
            
            -- lw
            when "100011" => 
                RegWrite <= '1';
                RegDst   <= '0';
                Branch   <= '0';
                MemRead  <= '1';
                MemtoReg <= '1';
                MemWrite <= '0';
                ALUSrc   <= '1';
                Jump     <= '0';
                ALUOp    <= "00"; -- ALUOp for lw/sw (add)
                
            -- sw 
            when "101011" => 
                RegWrite <= '0';
                RegDst   <= '0'; -- Typically 'X' or don't care, but setting to 0 is safe
                Branch   <= '0';
                MemRead  <= '0';
                MemtoReg <= '0'; -- Typically 'X'
                MemWrite <= '1';
                ALUSrc   <= '1';
                Jump     <= '0';
                ALUOp    <= "00"; -- ALUOp for lw/sw (add)

            -- beq 
            when "000100" => 
                RegWrite <= '0';
                RegDst   <= '0'; -- Typically 'X'
                Branch   <= '1';
                MemRead  <= '0';
                MemtoReg <= '0'; -- Typically 'X'
                MemWrite <= '0';
                ALUSrc   <= '0';
                Jump     <= '0';
                ALUOp    <= "01"; -- ALUOp for beq (subtract)
          
            -- jump
            when "000010" =>
                RegWrite <= '0';
                RegDst   <= '0'; -- Typically 'X'
                Branch   <= '0';
                MemRead  <= '0';
                MemtoReg <= '0'; -- Typically 'X'
                MemWrite <= '0';
                ALUSrc   <= '0'; -- Typically 'X'
                Jump     <= '1';
                ALUOp    <= "00"; -- ALUOp can be anything, ALU result not used for main path
		
            -- otros (other opcodes - default to safe/NOP-like values)
            when others =>		
                RegWrite <= '0';
                RegDst   <= '0';
                Branch   <= '0';
                MemRead  <= '0';
                MemtoReg <= '0';
                MemWrite <= '0';
                ALUSrc   <= '0';
                Jump     <= '0';
                ALUOp    <= "00"; -- Default ALUOp
        end case;
    end process;

    -- Assign the generated 2-bit ALUOp to the output port
    ALUOp_o <= ALUOp;

    -- The second process that generated the 4-bit ALUControl based on ALUOp and Funct is removed.
    -- That logic is now in the separate ALUControl module.

end architecture Behavioral;
